library ieee;
use ieee.std_logic_1164.all;

library unisim;
use unisim.vcomponents.all;

library unimacro;
use unimacro.vcomponents.all;


entity VgaCharacterRom is
    port (  clk : in std_logic;
            rst : in std_logic;
            char : in std_logic_vector(7 downto 0);
            pixelColumn : in std_logic_vector(2 downto 0);
            pixelRow : in std_logic_vector(3 downto 0);
            en : in std_logic;
            pixel : out std_logic);
end VgaCharacterRom;

architecture Structure of VgaCharacterRom is

signal address : std_logic_vector(14 downto 0);
signal pixel_vect : std_logic_vector(0 downto 0);

begin

    i_CharacterRom : BRAM_SINGLE_MACRO
        generic map (   BRAM_SIZE => "36Kb",
                        DEVICE => "7SERIES",
                        DO_REG => 0,
                        INIT => X"000000000000000000",
                        WRITE_WIDTH => 1,
                        READ_WIDTH => 1,
                        INIT_00 => X"000000007E818199BD8181A5817E000000000000000000000000000000000000",
                        INIT_01 => X"00000000081C3E7F7F7F7F3600000000000000007EFFFFE7C3FFFFDBFF7E0000",
                        INIT_02 => X"000000003C1818E7E7E73C3C180000000000000000081C3E7F3E1C0800000000",
                        INIT_03 => X"000000000000183C3C18000000000000000000003C18187EFFFF7E3C18000000",
                        INIT_04 => X"00000000003C664242663C0000000000FFFFFFFFFFFFE7C3C3E7FFFFFFFFFFFF",
                        INIT_05 => X"000000001E333333331E4C5870780000FFFFFFFFFFC399BDBD99C3FFFFFFFFFF",
                        INIT_06 => X"00000000070F0E0C0C0C0CFCCCFC00000000000018187E183C666666663C0000",
                        INIT_07 => X"000000001818DB3CE73CDB18180000000000000367E7E6C6C6C6C6FEC6FE0000",
                        INIT_08 => X"00000000406070787C7F7C7870604000000000000103070F1F7F1F0F07030100",
                        INIT_09 => X"000000006666006666666666666600000000000000183C7E1818187E3C180000",
                        INIT_0A => X"0000003E63301C366363361C06633E0000000000D8D8D8D8D8DEDBDBDBFE0000",
                        INIT_0B => X"000000007E183C7E1818187E3C180000000000007F7F7F7F0000000000000000",
                        INIT_0C => X"00000000183C7E18181818181818000000000000181818181818187E3C180000",
                        INIT_0D => X"0000000000000C067F060C000000000000000000000018307F30180000000000",
                        INIT_0E => X"00000000000014367F361400000000000000000000007F030303000000000000",
                        INIT_0F => X"0000000000081C1C3E3E7F7F0000000000000000007F7F3E3E1C1C0800000000",
                        INIT_10 => X"000000001818001818183C3C3C18000000000000000000000000000000000000",
                        INIT_11 => X"0000000036367F3636367F363600000000000000000000000000002466666600",
                        INIT_12 => X"000000006163060C1830634300000000000018183E636160603E0343633E1818",
                        INIT_13 => X"0000000000000000000000060C0C0C00000000006E3333333B6E1C36361C0000",
                        INIT_14 => X"000000000C18303030303030180C00000000000030180C0C0C0C0C0C18300000",
                        INIT_15 => X"00000000000018187E18180000000000000000000000663CFF3C660000000000",
                        INIT_16 => X"00000000000000007F000000000000000000000C181818000000000000000000",
                        INIT_17 => X"000000000103060C183060400000000000000000181800000000000000000000",
                        INIT_18 => X"000000007E1818181818181E1C180000000000001C3663636B6B6363361C0000",
                        INIT_19 => X"000000003E636060603C6060633E0000000000007F6303060C183060633E0000",
                        INIT_1A => X"000000003E636060603F0303037F000000000000783030307F33363C38300000",
                        INIT_1B => X"000000000C0C0C0C18306060637F0000000000003E636363633F0303061C0000",
                        INIT_1C => X"000000001E306060607E6363633E0000000000003E636363633E6363633E0000",
                        INIT_1D => X"000000000C181800000018180000000000000000001818000000181800000000",
                        INIT_1E => X"000000000000007E00007E0000000000000000006030180C060C183060000000",
                        INIT_1F => X"000000001818001818183063633E000000000000060C18306030180C06000000",
                        INIT_20 => X"00000000636363637F6363361C080000000000003E033B7B7B7B63633E000000",
                        INIT_21 => X"000000003C66430303030343663C0000000000003F666666663E6666663F0000",
                        INIT_22 => X"000000007F664606161E1646667F0000000000001F36666666666666361F0000",
                        INIT_23 => X"000000005C6663637B030343663C0000000000000F060606161E1646667F0000",
                        INIT_24 => X"000000003C18181818181818183C00000000000063636363637F636363630000",
                        INIT_25 => X"00000000676666361E1E366666670000000000001E3333333030303030780000",
                        INIT_26 => X"0000000063636363636B7F7F77630000000000007F66460606060606060F0000",
                        INIT_27 => X"000000003E63636363636363633E00000000000063636363737B7F6F67630000",
                        INIT_28 => X"000070303E7B6B6363636363633E0000000000000F060606063E6666663F0000",
                        INIT_29 => X"000000003E636360301C0663633E00000000000067666666363E6666663F0000",
                        INIT_2A => X"000000003E6363636363636363630000000000003C1818181818185A7E7E0000",
                        INIT_2B => X"0000000036777F6B6B6B63636363000000000000081C36636363636363630000",
                        INIT_2C => X"000000003C181818183C666666660000000000006363363E1C1C3E3663630000",
                        INIT_2D => X"000000003C0C0C0C0C0C0C0C0C3C0000000000007F6343060C183061637F0000",
                        INIT_2E => X"000000003C30303030303030303C000000000000406070381C0E070301000000",
                        INIT_2F => X"0000FF0000000000000000000000000000000000000000000000000063361C08",
                        INIT_30 => X"000000006E3333333E301E000000000000000000000000000000000000180C0C",
                        INIT_31 => X"000000003E63030303633E0000000000000000003E66666666361E0606070000",
                        INIT_32 => X"000000003E6303037F633E0000000000000000006E33333333363C3030380000",
                        INIT_33 => X"001E33303E33333333336E0000000000000000000F060606060F0626361C0000",
                        INIT_34 => X"000000003C18181818181C00181800000000000067666666666E360606070000",
                        INIT_35 => X"000000006766361E1E36660606070000003C6666606060606060700060600000",
                        INIT_36 => X"00000000636B6B6B6B7F370000000000000000003C18181818181818181C0000",
                        INIT_37 => X"000000003E63636363633E0000000000000000006666666666663B0000000000",
                        INIT_38 => X"007830303E33333333336E0000000000000F06063E66666666663B0000000000",
                        INIT_39 => X"000000003E63301C06633E0000000000000000000F060606666E3B0000000000",
                        INIT_3A => X"000000006E333333333333000000000000000000386C0C0C0C0C3F0C0C080000",
                        INIT_3B => X"00000000367F6B6B6B6363000000000000000000183C66666666660000000000",
                        INIT_3C => X"001F30607E63636363636300000000000000000063361C1C1C36630000000000",
                        INIT_3D => X"0000000070181818180E181818700000000000007F63060C18337F0000000000",
                        INIT_3E => X"000000000E18181818701818180E000000000000181818181800181818180000",
                        INIT_3F => X"00000000007F636363361C08000000000000000000000000000000003B6E0000",
                        INIT_40 => X"000000006E333333333333000033000000003E60303C664303030343663C0000",
                        INIT_41 => X"000000006E3333333E301E00361C0800000000003E6303037F633E000C183000",
                        INIT_42 => X"000000006E3333333E301E00180C0600000000006E3333333E301E0000330000",
                        INIT_43 => X"0000003C60303C660606663C00000000000000006E3333333E301E001C361C00",
                        INIT_44 => X"000000003E6303037F633E0000630000000000003E6303037F633E00361C0800",
                        INIT_45 => X"000000003C18181818181C0000660000000000003E6303037F633E00180C0600",
                        INIT_46 => X"000000003C18181818181C00180C0600000000003C18181818181C00663C1800",
                        INIT_47 => X"000000006363637F6363361C001C361C000000006363637F6363361C08006300",
                        INIT_48 => X"00000000761B1B7E6C6E330000000000000000007F6606063E06667F00060C18",
                        INIT_49 => X"000000003E63636363633E00361C08000000000073333333337F3333367C0000",
                        INIT_4A => X"000000003E63636363633E00180C0600000000003E63636363633E0000630000",
                        INIT_4B => X"000000006E33333333333300180C0600000000006E33333333333300331E0C00",
                        INIT_4C => X"000000003E636363636363633E006300001E30607E6363636363630000630000",
                        INIT_4D => X"0000000018183C66060606663C181800000000003E6363636363636363006300",
                        INIT_4E => X"000000001818187E187E183C66660000000000003F67060606060F0626361C00",
                        INIT_4F => X"00000E1B18181818187E181818D8700000000000633333337B33231F33331F00",
                        INIT_50 => X"000000003C18181818181C000C183000000000006E3333333E301E00060C1800",
                        INIT_51 => X"000000006E33333333333300060C1800000000003E63636363633E00060C1800",
                        INIT_52 => X"00000000636363737B7F6F6763003B6E000000006666666666663B003B6E0000",
                        INIT_53 => X"0000000000000000003E001C36361C000000000000000000007E007C36363C00",
                        INIT_54 => X"0000000000030303037F000000000000000000003E636303060C0C000C0C0000",
                        INIT_55 => X"00007C1830613B060C183363430303000000000000606060607F000000000000",
                        INIT_56 => X"00000000183C3C3C1818180018180000000060607C7973660C18336343030300",
                        INIT_57 => X"0000000000001B366C361B00000000000000000000006C361B366C0000000000",
                        INIT_58 => X"55AA55AA55AA55AA55AA55AA55AA55AA22882288228822882288228822882288",
                        INIT_59 => X"18181818181818181818181818181818EEBBEEBBEEBBEEBBEEBBEEBBEEBBEEBB",
                        INIT_5A => X"18181818181818181F181F181818181818181818181818181F18181818181818",
                        INIT_5B => X"6C6C6C6C6C6C6C6C7F000000000000006C6C6C6C6C6C6C6C6F6C6C6C6C6C6C6C",
                        INIT_5C => X"6C6C6C6C6C6C6C6C6F606F6C6C6C6C6C18181818181818181F181F0000000000",
                        INIT_5D => X"6C6C6C6C6C6C6C6C6F607F00000000006C6C6C6C6C6C6C6C6C6C6C6C6C6C6C6C",
                        INIT_5E => X"00000000000000007F6C6C6C6C6C6C6C00000000000000007F606F6C6C6C6C6C",
                        INIT_5F => X"18181818181818181F0000000000000000000000000000001F181F1818181818",
                        INIT_60 => X"0000000000000000FF181818181818180000000000000000F818181818181818",
                        INIT_61 => X"1818181818181818F8181818181818181818181818181818FF00000000000000",
                        INIT_62 => X"1818181818181818FF181818181818180000000000000000FF00000000000000",
                        INIT_63 => X"6C6C6C6C6C6C6C6CEC6C6C6C6C6C6C6C1818181818181818F818F81818181818",
                        INIT_64 => X"6C6C6C6C6C6C6C6CEC0CFC00000000000000000000000000FC0CEC6C6C6C6C6C",
                        INIT_65 => X"6C6C6C6C6C6C6C6CEF00FF00000000000000000000000000FF00EF6C6C6C6C6C",
                        INIT_66 => X"0000000000000000FF00FF00000000006C6C6C6C6C6C6C6CEC0CEC6C6C6C6C6C",
                        INIT_67 => X"0000000000000000FF00FF18181818186C6C6C6C6C6C6C6CEF00EF6C6C6C6C6C",
                        INIT_68 => X"1818181818181818FF00FF00000000000000000000000000FF6C6C6C6C6C6C6C",
                        INIT_69 => X"0000000000000000FC6C6C6C6C6C6C6C6C6C6C6C6C6C6C6CFF00000000000000",
                        INIT_6A => X"1818181818181818F818F800000000000000000000000000F818F81818181818",
                        INIT_6B => X"6C6C6C6C6C6C6C6CFF6C6C6C6C6C6C6C6C6C6C6C6C6C6C6CFC00000000000000",
                        INIT_6C => X"00000000000000001F181818181818181818181818181818FF18FF1818181818",
                        INIT_6D => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1818181818181818F800000000000000",
                        INIT_6E => X"0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0FFFFFFFFFFFFFFFFFFF00000000000000",
                        INIT_6F => X"000000000000000000FFFFFFFFFFFFFFF0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0",
                        INIT_70 => X"0000000033636363331B3333331E0000000000006E3B1B1B1B3B6E0000000000",
                        INIT_71 => X"00000000363636363636367F00000000000000000303030303030363637F0000",
                        INIT_72 => X"000000000E1B1B1B1B1B7E0000000000000000007F63060C180C06637F000000",
                        INIT_73 => X"000000001818181818183B6E000000000000000306063E666666666600000000",
                        INIT_74 => X"000000001C3663637F6363361C000000000000007E183C6666663C187E000000",
                        INIT_75 => X"000000003C666666667C30180C780000000000007736363636636363361C0000",
                        INIT_76 => X"0000000003067ECFDBDB7E60C00000000000000000007EDBDBDB7E0000000000",
                        INIT_77 => X"0000000063636363636363633E00000000000000380C0606063E06060C380000",
                        INIT_78 => X"00000000FF000018187E18180000000000000000007F00007F00007F00000000",
                        INIT_79 => X"000000007E0030180C060C1830000000000000007E000C18306030180C000000",
                        INIT_7A => X"000000000E1B1B1B18181818181818181818181818181818181818D8D8700000",
                        INIT_7B => X"0000000000003B6E003B6E000000000000000000001818007E00181800000000",
                        INIT_7C => X"0000000000000018180000000000000000000000000000000000001C36361C00",
                        INIT_7D => X"00000000383C3636373030303030F00000000000000000180000000000000000",
                        INIT_7E => X"0000000000000000001F13060C1B0E0000000000000000000036363636361B00",
                        INIT_7F => X"0000000000000000000000000000000000000000003E3E3E3E3E3E3E00000000")
        port map (  CLK => clk,
                    RST => '0',
                    DO => pixel_vect,
                    ADDR => address,
                    EN => en,
                    REGCE => '0',
                    DI => "0",
                    WE => "0");

    address <= char & pixelRow & pixelColumn;
    pixel <= pixel_vect(0);

end Structure;
